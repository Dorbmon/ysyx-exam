`include "vsrc/template.v"

module ysyx_22041207_top (
  input [31:0] inst,
  output reg [31:0] pc
);
endmodule