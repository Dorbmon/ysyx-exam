module ysyx_22041207_auipc(
    input is
);

endmodule